# ========== APP ==========
APP_TITLE="Mordzix PRO ULTRA"
APP_VERSION=3.2.0
ALLOWED_ORIGINS=*

# ========== AUTH ==========
AUTH_TOKEN=ssjjMijaja6969

# ========== LOGGING / DEBUG ==========
LOGLEVEL=INFO
IMG_DEBUG=0
PSY_DEBUG=0

# ========== CORE PATHS ==========
OUT_DIR=/workspace/mrd69/overmind/output
WRITER_OUT_DIR=/workspace/mrd69/overmind/output/writing
IMG_OUT_DIR=/workspace/mrd69/overmind/output/images
MEM_DIR=/workspace/mrd69/overmind/memory
LTM_DB_PATH=/workspace/mrd69/overmind/memory/ltm.db
PROMPT_BASE_RULES=/workspace/mrd69/overmind/prompts/mordzix_system.txt

# ========== DEV TOOL (programista.py) ==========
DEV_OUT_DIR=/workspace/mrd69/overmind/output/dev
DEV_SAVE_JSON=1
DEV_ZIP_EXPORT=1
DEV_MAX_WORKERS=8
DEV_TOOL_TIMEOUT=18
DEV_FAIL_MI=0

# ========== LLM (MAIN – DeepInfra/OpenAI compatible) ==========
export 
LLM_BASE_URL=https://api.deepinfra.com/v1/openai 
LLM_HTTP_TIMEOUT_S=60 LLM_TIMEOUT=60 
LLM_RETRIES=3 LLM_BACKOFF_S=2 LLM_MAX_CONC=4 
LLM_CACHE_TTL_S=300 LLM_COST_PROMPT_PER_1K=0 
LLM_COST_COMP_PER_1K=0 LLM_JOURNAL=0 export 
LLM_MODEL=Qwen/Qwen2.5-72B-Instruct export 
LLM_API_KEY=aMT2CsbRlkpqU9ZaoIPgTvrL4pa7pM8H# 
Embeddings 
LLM_EMBED_URL=https://api.openai.com/v1/embeddings 
LLM_EMBED_MODEL=text-embedding-3-large

# Reranker
LLM_RERANK_URL=https://api.deepinfra.com/v1/rerank
LLM_RERANK_KEY=nkQfwzC0zwjglJpwgbo3SQIfpTZIfv2u

# ========== MINI LLM (BG tasks – Qwen 4B) ==========
MINI_LLM_BASE_URL=https://api.deepinfra.com/v1/openai
MINI_LLM_API_KEY=nkQfwzC0zwjglJpwgbo3SQIfpTZIfv2u
MINI_LLM_MODEL=Qwen/Qwen2.5-4B-Instruct
MINI_LLM_TIMEOUT_S=30
MINI_LLM_RETRIES=2
MINI_LLM_BACKOFF_S=1
USE_MINI_FOR_BG=1

# ========== OpenAI (fallback) ==========
OPENAI_BASE_URL=https://api.openai.com/v1
OPENAI_API_KEY=sk-proj-EmKhjmI2SHrDjK75ocjI5OuKI_Uea7qQO-d7t0
OPENAI_KEY=sk-proj-EmKhjmI2SHrDjK75ocjI5OuKI_Uea7qQO-d7t0

# ========== Google / Vertex / Gemini ==========
GOOGLE_API_KEY=AIzaSyA01GWKXRX9x_MyRnoBUwCvFqnjwZa-Bao
GOOGLE_BOOKS_KEY=AlzaSyC8vsWs3XzfNWrU1gQNNk2QwZQYKCFS3Es
GOOGLE_CSE_KEY=
GOOGLE_CSE_CX=
GOOGLE_CLOUD_PROJECT=
GOOGLE_CLOUD_LOCATION=
GOOGLE_CLOUD_STORAGE_BUCKET=
GOOGLE_CLOUD_BQ_DATASET=
GOOGLE_OAUTH_TOKEN=
GOOGLE_GENAI_MODEL=
GOOGLE_GENAI_USE_VERTEXAI=
GOOGLE_GENAI_FOMC_AGENT_LOG_LEVEL=
GOOGLE_GENAI_FOMC_AGENT_TIMESERIES_CODES=

# Gemini (API bez Vertex) – jeśli używasz:
GEMINI_API_KEY=
GEMINI_MODEL=
GEMINI_EMBED_MODEL=

# Vertex AI (jeśli używasz):
VERTEX_GEMINI_KEY=AlzaSyAKouyWh_tQ2LppvU54DJF97KpzgHHjYCA
VERTEX_MODEL=
VERTEX_PROJECT=
VERTEX_LOCATION=
VERTEX_TOKEN=
VERTEX_OAUTH_BEARER=

# ========== Web / RAG / Crawling ==========
WEB_USER_AGENT="MordzixBot/1.0"
WEB_HTTP_TIMEOUT=45
HTTP_TIMEOUT=60
TIMEOUT_HTTP=60
AUTO_FETCH=
AUTO_MAX_CHARS=
AUTO_MIN_CHARS=
AUTO_TOPK=
AUTO_TAGS=
CACHE_TTL=
RAG_TOPK=5
RAG_CACHE_TTL_MIN=30
RAG_PAR_SCRAPE=1
DISABLE_WEB_DRIVER=

SERPAPI_KEY=a5cb3592980e0ff9042a0be2d3f7df2768bd93913252
FIRECRAWL_KEY=fc-ec025f3a447c6878bee6926b49c17d3

# ========== Maps / Travel / Weather ==========
OVERPASS_URL=https://overpass-api.de/api/interpreter
GOOGLE_PLACES_API_KEY=
GOOGLE_PLACES_KEY=
MAPS_STATIC_KEY=AlzaSyCvwN2RWhEJ2t2JHZQQQztoaDZHpFS6Pgl
MAPTILER_KEY=wczEnYV9dtQUGgduQIxPoAQDp2wH4qehTPQuL
TRAVEL_PARTNER_KEY=AlzaSyCbpKUI1Vt9sGmmU0eRhgLpUtevegXWgy8

TRAVEL_CACHE_TTL_MIN=120
TRAVEL_MAX_RESULTS=
TRAVEL_NEARBY_RADIUS=
TRAVEL_CONCIERGE_SCENARIO=
TRAVEL_FOOD_PREFS=ramen,pizza,tapas,vegan,seafood
TRAVEL_HOTEL_PREFS=marriott,hilton,ibis,aparthotel,hostel

OPENWEATHER_KEY=cbe8e0a228ba0697f1cf5cd64bbef3e6
VISUAL_CROSSING_KEY=MHSNYKTD26EDJVPWZ3SM5HAG9

# ========== Graphics (Stability + HF) ==========
STABILITY_API_KEY=sk-WslJMSme2LXkvXI8B7660lCfsTQt9VPxdRA4JovF
STABILITY_KEY=sk-WslJMSme2LXkvXI8B7660lCfsTQt9VPxdRA4JovF
STABILITY_ENGINE=stable-diffusion-xl-1024-v1-0
STABILITY_SD3_ENDPOINT=

HF_TOKEN=hf_VTyPVDyhszhoEhIZApLQTxQBCishBbZC1T
HUGGINGFACE_API_KEY=hf_VTyPVDyhszhoEhIZApLQTxQBCishBbZC1T
HF_TXT2IMG_MODEL=
HF_IMG2IMG_MODEL=
HF_INPAINT_MODEL=
HF_OUTPAINT_MODEL=
HF_CONTROLNET_MODEL=
HF_DEPTH_MODEL=

IMG_PREVIEW_W=768
IMG_TOPN=4

# ========== Crypto / Finance ==========
COINGECKO_VS=
PORTFOLIO_USD=
RISK_CAP_PCT=
ETHERSCAN_API_KEY=Q86S7ZHDKQRXUGMAQIX21YUA7TXE4SFZ9V
WHALE_ADDRS=

# ========== OSS / Code Quality ==========
OSS_INDEX_TOKEN=3f476a939384bfc0db197e368c3e4588a98d2019
SONAR_TOKEN=44e5f20fc65ccd66c5a65a7d8b133867bbb88f02

# ========== Telegram / Notyfikacje ==========
TELEGRAM_BOT_TOKEN=
TELEGRAM_CHAT_ID=
SERVE_WEB_INTERFACE=

# ========== Memory / Psychika ==========
MEM_NS=default
MEM_STM_WINDOW=16
MEM_LTM_MAX=2000
LTM_MIN_CONF=0.35
LTM_DB_MAX_BYTES=104857600

PSY_ENCRYPT_KEY=dev_psy_key_change_me
PSY_BANDIT=
PSY_BRIDGE_FETCH=
PSY_BRIDGE_MODE=
PSY_BRIDGE_TOPK=
PSY_COMPASSION=
PSY_DUTY=
PSY_EXPLORATION=
PSY_GOAL_WEIGHT=
PSY_HONOR=
PSY_MAX_OPTIONS=
PSY_MORALITY=
PSY_PARETO=
PSY_PRESET=
PSY_PRIDE=
PSY_RECIPROCITY=
PSY_REGRET=
PSY_RELIEF=
PSY_RISK_AVERSION=
PSY_SEED=
PSY_UNWRAP=
PSY_WEB_WHITELIST=

STM_KEEP_TAIL=6
STM_MAX_TURNS=16
HISTORY_MAX_TURNS=32
MAX_EP_LINES=
MAX_ITERATIONS=
MAX_LTM_FACTS=

# ========== Analytics / Agents / Models ==========
ANALYTICS_AGENT_MODEL=
ROOT_AGENT_MODEL=
AGENT_ENGINE_ID=
GENAI_MODEL=
MODEL=
SCORE_THRESHOLD=

# ========== Data / BigQuery / Dataform (jeśli używasz) ==========
GCP_PROJECT_ID=
BQ_DATA_PROJECT_ID=
BQ_COMPUTE_PROJECT_ID=
BQ_DATASET_ID=
DATASET_ID=
TABLE_ID=
GOOGLE_CLOUD_BQ_DATASET=
DATAFORM_REPOSITORY_NAME=
DATAFORM_WORKSPACE_NAME=
BQML_AGENT_MODEL=
BQML_RAG_CORPUS_NAME=
BASELINE_NL2SQL_MODEL=
CHASE_NL2SQL_MODEL=
NL2SQL_METHOD=

# ========== Dedup / Rerank / Search heur ==========
DEDUP_EMB=
DEDUP_EMB_THR=
DEDUP_TFIDF=
DEDUP_TFIDF_THR=
DEDUP_NORM_HASH=
HYBRID_MODE=
HYBRID_W_WEB=
HYBRID_W_MEM=
HYBRID_W_HEUR=
RECALL_TOPK_PER_SRC=

# ========== Misc Tools / OCR / Images ==========
OCR_LANG=
IMG_HTTP_TIMEOUT=30

# ========== Background worker ==========
BG_AUTOSTART=1
BG_QUEUE_DIR=/workspace/mrd69/overmind/queue

# ========== Optional Keys, które podałeś (aliasy) ==========
BOOKS_API_KEY=AlzaSyC8vsWs3XzfNWrU1gQNNk2QwZQYKCFS3Es
MAPS_STATIC_API_KEY=AlzaSyCvwN2RWhEJ2t2JHZQQQztoaDZHpFS6Pgl
GENERATIVE_LANGUAGE_API_KEY=AIzaSyA01GWKXRX9x_MyRnoBUwCvFqnjwZa-Bao
TRAVEL_PARTNER_API_KEY=AlzaSyCbpKUI1Vt9sGmmU0eRhgLpUtevegXWgy8

# ========== Not used / legacy toggles (zostaw puste jeśli niepotrzebne) ==========
ESRGAN_ON=
GFPGAN_ON=
IMAGEN_MODEL=
ADK_WHL_FILE=
CG_BASE=
CG_PAUSE=
CG_TIMEOUT=
CODE_INTERPRETER_EXTENSION_NAME=
DISABLE_WEB_DRIVER=
ERC20_CONTRACT=
GITHUB_PERSONAL_ACCESS_TOKEN=
IMG_SELFTEST_OUTDIR=
IMG_SELFTEST_PROMPT=
MCP_TOOLBOX_URL=
STAGING_BUCKET=
SESSION_SERVICE_URI=
SERVE_WEB_INTERFACE=
VAR=
WATCHLIST=
WEB_HTTP_TIMEOUT=
